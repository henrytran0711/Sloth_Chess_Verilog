module serializer(clk, in, load, w_en, data_out, move_counter_out,done);

  input clk;
  input [24191:0] in;
  input load;
  input w_en;
  output reg [31:0] data_out;
  output reg done;
  output reg [9:0] move_counter_out;
  reg [31:0] mem [755:0];
  reg [9:0] r_addr;
  reg [9:0] move_counter;
  
  initial begin
	 move_counter = 10'd000;
	 done = 1'b0;
	 
  end
  always @(posedge clk) begin
    if(load) begin
      r_addr = 10'b00000_00000;
      mem[10'd0] <= in[24191:24160];
      mem[10'd1] <= in[24159:24128];
      mem[10'd2] <= in[24127:24096];
      mem[10'd3] <= in[24095:24064];
      mem[10'd4] <= in[24063:24032];
      mem[10'd5] <= in[24031:24000];
      mem[10'd6] <= in[23999:23968];
      mem[10'd7] <= in[23967:23936];
      mem[10'd8] <= in[23935:23904];
      mem[10'd9] <= in[23903:23872];
      mem[10'd10] <= in[23871:23840];
      mem[10'd11] <= in[23839:23808];
      mem[10'd12] <= in[23807:23776];
      mem[10'd13] <= in[23775:23744];
      mem[10'd14] <= in[23743:23712];
      mem[10'd15] <= in[23711:23680];
      mem[10'd16] <= in[23679:23648];
      mem[10'd17] <= in[23647:23616];
      mem[10'd18] <= in[23615:23584];
      mem[10'd19] <= in[23583:23552];
      mem[10'd20] <= in[23551:23520];
      mem[10'd21] <= in[23519:23488];
      mem[10'd22] <= in[23487:23456];
      mem[10'd23] <= in[23455:23424];
      mem[10'd24] <= in[23423:23392];
      mem[10'd25] <= in[23391:23360];
      mem[10'd26] <= in[23359:23328];
      mem[10'd27] <= in[23327:23296];
      mem[10'd28] <= in[23295:23264];
      mem[10'd29] <= in[23263:23232];
      mem[10'd30] <= in[23231:23200];
      mem[10'd31] <= in[23199:23168];
      mem[10'd32] <= in[23167:23136];
      mem[10'd33] <= in[23135:23104];
      mem[10'd34] <= in[23103:23072];
      mem[10'd35] <= in[23071:23040];
      mem[10'd36] <= in[23039:23008];
      mem[10'd37] <= in[23007:22976];
      mem[10'd38] <= in[22975:22944];
      mem[10'd39] <= in[22943:22912];
      mem[10'd40] <= in[22911:22880];
      mem[10'd41] <= in[22879:22848];
      mem[10'd42] <= in[22847:22816];
      mem[10'd43] <= in[22815:22784];
      mem[10'd44] <= in[22783:22752];
      mem[10'd45] <= in[22751:22720];
      mem[10'd46] <= in[22719:22688];
      mem[10'd47] <= in[22687:22656];
      mem[10'd48] <= in[22655:22624];
      mem[10'd49] <= in[22623:22592];
      mem[10'd50] <= in[22591:22560];
      mem[10'd51] <= in[22559:22528];
      mem[10'd52] <= in[22527:22496];
      mem[10'd53] <= in[22495:22464];
      mem[10'd54] <= in[22463:22432];
      mem[10'd55] <= in[22431:22400];
      mem[10'd56] <= in[22399:22368];
      mem[10'd57] <= in[22367:22336];
      mem[10'd58] <= in[22335:22304];
      mem[10'd59] <= in[22303:22272];
      mem[10'd60] <= in[22271:22240];
      mem[10'd61] <= in[22239:22208];
      mem[10'd62] <= in[22207:22176];
      mem[10'd63] <= in[22175:22144];
      mem[10'd64] <= in[22143:22112];
      mem[10'd65] <= in[22111:22080];
      mem[10'd66] <= in[22079:22048];
      mem[10'd67] <= in[22047:22016];
      mem[10'd68] <= in[22015:21984];
      mem[10'd69] <= in[21983:21952];
      mem[10'd70] <= in[21951:21920];
      mem[10'd71] <= in[21919:21888];
      mem[10'd72] <= in[21887:21856];
      mem[10'd73] <= in[21855:21824];
      mem[10'd74] <= in[21823:21792];
      mem[10'd75] <= in[21791:21760];
      mem[10'd76] <= in[21759:21728];
      mem[10'd77] <= in[21727:21696];
      mem[10'd78] <= in[21695:21664];
      mem[10'd79] <= in[21663:21632];
      mem[10'd80] <= in[21631:21600];
      mem[10'd81] <= in[21599:21568];
      mem[10'd82] <= in[21567:21536];
      mem[10'd83] <= in[21535:21504];
      mem[10'd84] <= in[21503:21472];
      mem[10'd85] <= in[21471:21440];
      mem[10'd86] <= in[21439:21408];
      mem[10'd87] <= in[21407:21376];
      mem[10'd88] <= in[21375:21344];
      mem[10'd89] <= in[21343:21312];
      mem[10'd90] <= in[21311:21280];
      mem[10'd91] <= in[21279:21248];
      mem[10'd92] <= in[21247:21216];
      mem[10'd93] <= in[21215:21184];
      mem[10'd94] <= in[21183:21152];
      mem[10'd95] <= in[21151:21120];
      mem[10'd96] <= in[21119:21088];
      mem[10'd97] <= in[21087:21056];
      mem[10'd98] <= in[21055:21024];
      mem[10'd99] <= in[21023:20992];
      mem[10'd100] <= in[20991:20960];
      mem[10'd101] <= in[20959:20928];
      mem[10'd102] <= in[20927:20896];
      mem[10'd103] <= in[20895:20864];
      mem[10'd104] <= in[20863:20832];
      mem[10'd105] <= in[20831:20800];
      mem[10'd106] <= in[20799:20768];
      mem[10'd107] <= in[20767:20736];
      mem[10'd108] <= in[20735:20704];
      mem[10'd109] <= in[20703:20672];
      mem[10'd110] <= in[20671:20640];
      mem[10'd111] <= in[20639:20608];
      mem[10'd112] <= in[20607:20576];
      mem[10'd113] <= in[20575:20544];
      mem[10'd114] <= in[20543:20512];
      mem[10'd115] <= in[20511:20480];
      mem[10'd116] <= in[20479:20448];
      mem[10'd117] <= in[20447:20416];
      mem[10'd118] <= in[20415:20384];
      mem[10'd119] <= in[20383:20352];
      mem[10'd120] <= in[20351:20320];
      mem[10'd121] <= in[20319:20288];
      mem[10'd122] <= in[20287:20256];
      mem[10'd123] <= in[20255:20224];
      mem[10'd124] <= in[20223:20192];
      mem[10'd125] <= in[20191:20160];
      mem[10'd126] <= in[20159:20128];
      mem[10'd127] <= in[20127:20096];
      mem[10'd128] <= in[20095:20064];
      mem[10'd129] <= in[20063:20032];
      mem[10'd130] <= in[20031:20000];
      mem[10'd131] <= in[19999:19968];
      mem[10'd132] <= in[19967:19936];
      mem[10'd133] <= in[19935:19904];
      mem[10'd134] <= in[19903:19872];
      mem[10'd135] <= in[19871:19840];
      mem[10'd136] <= in[19839:19808];
      mem[10'd137] <= in[19807:19776];
      mem[10'd138] <= in[19775:19744];
      mem[10'd139] <= in[19743:19712];
      mem[10'd140] <= in[19711:19680];
      mem[10'd141] <= in[19679:19648];
      mem[10'd142] <= in[19647:19616];
      mem[10'd143] <= in[19615:19584];
      mem[10'd144] <= in[19583:19552];
      mem[10'd145] <= in[19551:19520];
      mem[10'd146] <= in[19519:19488];
      mem[10'd147] <= in[19487:19456];
      mem[10'd148] <= in[19455:19424];
      mem[10'd149] <= in[19423:19392];
      mem[10'd150] <= in[19391:19360];
      mem[10'd151] <= in[19359:19328];
      mem[10'd152] <= in[19327:19296];
      mem[10'd153] <= in[19295:19264];
      mem[10'd154] <= in[19263:19232];
      mem[10'd155] <= in[19231:19200];
      mem[10'd156] <= in[19199:19168];
      mem[10'd157] <= in[19167:19136];
      mem[10'd158] <= in[19135:19104];
      mem[10'd159] <= in[19103:19072];
      mem[10'd160] <= in[19071:19040];
      mem[10'd161] <= in[19039:19008];
      mem[10'd162] <= in[19007:18976];
      mem[10'd163] <= in[18975:18944];
      mem[10'd164] <= in[18943:18912];
      mem[10'd165] <= in[18911:18880];
      mem[10'd166] <= in[18879:18848];
      mem[10'd167] <= in[18847:18816];
      mem[10'd168] <= in[18815:18784];
      mem[10'd169] <= in[18783:18752];
      mem[10'd170] <= in[18751:18720];
      mem[10'd171] <= in[18719:18688];
      mem[10'd172] <= in[18687:18656];
      mem[10'd173] <= in[18655:18624];
      mem[10'd174] <= in[18623:18592];
      mem[10'd175] <= in[18591:18560];
      mem[10'd176] <= in[18559:18528];
      mem[10'd177] <= in[18527:18496];
      mem[10'd178] <= in[18495:18464];
      mem[10'd179] <= in[18463:18432];
      mem[10'd180] <= in[18431:18400];
      mem[10'd181] <= in[18399:18368];
      mem[10'd182] <= in[18367:18336];
      mem[10'd183] <= in[18335:18304];
      mem[10'd184] <= in[18303:18272];
      mem[10'd185] <= in[18271:18240];
      mem[10'd186] <= in[18239:18208];
      mem[10'd187] <= in[18207:18176];
      mem[10'd188] <= in[18175:18144];
      mem[10'd189] <= in[18143:18112];
      mem[10'd190] <= in[18111:18080];
      mem[10'd191] <= in[18079:18048];
      mem[10'd192] <= in[18047:18016];
      mem[10'd193] <= in[18015:17984];
      mem[10'd194] <= in[17983:17952];
      mem[10'd195] <= in[17951:17920];
      mem[10'd196] <= in[17919:17888];
      mem[10'd197] <= in[17887:17856];
      mem[10'd198] <= in[17855:17824];
      mem[10'd199] <= in[17823:17792];
      mem[10'd200] <= in[17791:17760];
      mem[10'd201] <= in[17759:17728];
      mem[10'd202] <= in[17727:17696];
      mem[10'd203] <= in[17695:17664];
      mem[10'd204] <= in[17663:17632];
      mem[10'd205] <= in[17631:17600];
      mem[10'd206] <= in[17599:17568];
      mem[10'd207] <= in[17567:17536];
      mem[10'd208] <= in[17535:17504];
      mem[10'd209] <= in[17503:17472];
      mem[10'd210] <= in[17471:17440];
      mem[10'd211] <= in[17439:17408];
      mem[10'd212] <= in[17407:17376];
      mem[10'd213] <= in[17375:17344];
      mem[10'd214] <= in[17343:17312];
      mem[10'd215] <= in[17311:17280];
      mem[10'd216] <= in[17279:17248];
      mem[10'd217] <= in[17247:17216];
      mem[10'd218] <= in[17215:17184];
      mem[10'd219] <= in[17183:17152];
      mem[10'd220] <= in[17151:17120];
      mem[10'd221] <= in[17119:17088];
      mem[10'd222] <= in[17087:17056];
      mem[10'd223] <= in[17055:17024];
      mem[10'd224] <= in[17023:16992];
      mem[10'd225] <= in[16991:16960];
      mem[10'd226] <= in[16959:16928];
      mem[10'd227] <= in[16927:16896];
      mem[10'd228] <= in[16895:16864];
      mem[10'd229] <= in[16863:16832];
      mem[10'd230] <= in[16831:16800];
      mem[10'd231] <= in[16799:16768];
      mem[10'd232] <= in[16767:16736];
      mem[10'd233] <= in[16735:16704];
      mem[10'd234] <= in[16703:16672];
      mem[10'd235] <= in[16671:16640];
      mem[10'd236] <= in[16639:16608];
      mem[10'd237] <= in[16607:16576];
      mem[10'd238] <= in[16575:16544];
      mem[10'd239] <= in[16543:16512];
      mem[10'd240] <= in[16511:16480];
      mem[10'd241] <= in[16479:16448];
      mem[10'd242] <= in[16447:16416];
      mem[10'd243] <= in[16415:16384];
      mem[10'd244] <= in[16383:16352];
      mem[10'd245] <= in[16351:16320];
      mem[10'd246] <= in[16319:16288];
      mem[10'd247] <= in[16287:16256];
      mem[10'd248] <= in[16255:16224];
      mem[10'd249] <= in[16223:16192];
      mem[10'd250] <= in[16191:16160];
      mem[10'd251] <= in[16159:16128];
      mem[10'd252] <= in[16127:16096];
      mem[10'd253] <= in[16095:16064];
      mem[10'd254] <= in[16063:16032];
      mem[10'd255] <= in[16031:16000];
      mem[10'd256] <= in[15999:15968];
      mem[10'd257] <= in[15967:15936];
      mem[10'd258] <= in[15935:15904];
      mem[10'd259] <= in[15903:15872];
      mem[10'd260] <= in[15871:15840];
      mem[10'd261] <= in[15839:15808];
      mem[10'd262] <= in[15807:15776];
      mem[10'd263] <= in[15775:15744];
      mem[10'd264] <= in[15743:15712];
      mem[10'd265] <= in[15711:15680];
      mem[10'd266] <= in[15679:15648];
      mem[10'd267] <= in[15647:15616];
      mem[10'd268] <= in[15615:15584];
      mem[10'd269] <= in[15583:15552];
      mem[10'd270] <= in[15551:15520];
      mem[10'd271] <= in[15519:15488];
      mem[10'd272] <= in[15487:15456];
      mem[10'd273] <= in[15455:15424];
      mem[10'd274] <= in[15423:15392];
      mem[10'd275] <= in[15391:15360];
      mem[10'd276] <= in[15359:15328];
      mem[10'd277] <= in[15327:15296];
      mem[10'd278] <= in[15295:15264];
      mem[10'd279] <= in[15263:15232];
      mem[10'd280] <= in[15231:15200];
      mem[10'd281] <= in[15199:15168];
      mem[10'd282] <= in[15167:15136];
      mem[10'd283] <= in[15135:15104];
      mem[10'd284] <= in[15103:15072];
      mem[10'd285] <= in[15071:15040];
      mem[10'd286] <= in[15039:15008];
      mem[10'd287] <= in[15007:14976];
      mem[10'd288] <= in[14975:14944];
      mem[10'd289] <= in[14943:14912];
      mem[10'd290] <= in[14911:14880];
      mem[10'd291] <= in[14879:14848];
      mem[10'd292] <= in[14847:14816];
      mem[10'd293] <= in[14815:14784];
      mem[10'd294] <= in[14783:14752];
      mem[10'd295] <= in[14751:14720];
      mem[10'd296] <= in[14719:14688];
      mem[10'd297] <= in[14687:14656];
      mem[10'd298] <= in[14655:14624];
      mem[10'd299] <= in[14623:14592];
      mem[10'd300] <= in[14591:14560];
      mem[10'd301] <= in[14559:14528];
      mem[10'd302] <= in[14527:14496];
      mem[10'd303] <= in[14495:14464];
      mem[10'd304] <= in[14463:14432];
      mem[10'd305] <= in[14431:14400];
      mem[10'd306] <= in[14399:14368];
      mem[10'd307] <= in[14367:14336];
      mem[10'd308] <= in[14335:14304];
      mem[10'd309] <= in[14303:14272];
      mem[10'd310] <= in[14271:14240];
      mem[10'd311] <= in[14239:14208];
      mem[10'd312] <= in[14207:14176];
      mem[10'd313] <= in[14175:14144];
      mem[10'd314] <= in[14143:14112];
      mem[10'd315] <= in[14111:14080];
      mem[10'd316] <= in[14079:14048];
      mem[10'd317] <= in[14047:14016];
      mem[10'd318] <= in[14015:13984];
      mem[10'd319] <= in[13983:13952];
      mem[10'd320] <= in[13951:13920];
      mem[10'd321] <= in[13919:13888];
      mem[10'd322] <= in[13887:13856];
      mem[10'd323] <= in[13855:13824];
      mem[10'd324] <= in[13823:13792];
      mem[10'd325] <= in[13791:13760];
      mem[10'd326] <= in[13759:13728];
      mem[10'd327] <= in[13727:13696];
      mem[10'd328] <= in[13695:13664];
      mem[10'd329] <= in[13663:13632];
      mem[10'd330] <= in[13631:13600];
      mem[10'd331] <= in[13599:13568];
      mem[10'd332] <= in[13567:13536];
      mem[10'd333] <= in[13535:13504];
      mem[10'd334] <= in[13503:13472];
      mem[10'd335] <= in[13471:13440];
      mem[10'd336] <= in[13439:13408];
      mem[10'd337] <= in[13407:13376];
      mem[10'd338] <= in[13375:13344];
      mem[10'd339] <= in[13343:13312];
      mem[10'd340] <= in[13311:13280];
      mem[10'd341] <= in[13279:13248];
      mem[10'd342] <= in[13247:13216];
      mem[10'd343] <= in[13215:13184];
      mem[10'd344] <= in[13183:13152];
      mem[10'd345] <= in[13151:13120];
      mem[10'd346] <= in[13119:13088];
      mem[10'd347] <= in[13087:13056];
      mem[10'd348] <= in[13055:13024];
      mem[10'd349] <= in[13023:12992];
      mem[10'd350] <= in[12991:12960];
      mem[10'd351] <= in[12959:12928];
      mem[10'd352] <= in[12927:12896];
      mem[10'd353] <= in[12895:12864];
      mem[10'd354] <= in[12863:12832];
      mem[10'd355] <= in[12831:12800];
      mem[10'd356] <= in[12799:12768];
      mem[10'd357] <= in[12767:12736];
      mem[10'd358] <= in[12735:12704];
      mem[10'd359] <= in[12703:12672];
      mem[10'd360] <= in[12671:12640];
      mem[10'd361] <= in[12639:12608];
      mem[10'd362] <= in[12607:12576];
      mem[10'd363] <= in[12575:12544];
      mem[10'd364] <= in[12543:12512];
      mem[10'd365] <= in[12511:12480];
      mem[10'd366] <= in[12479:12448];
      mem[10'd367] <= in[12447:12416];
      mem[10'd368] <= in[12415:12384];
      mem[10'd369] <= in[12383:12352];
      mem[10'd370] <= in[12351:12320];
      mem[10'd371] <= in[12319:12288];
      mem[10'd372] <= in[12287:12256];
      mem[10'd373] <= in[12255:12224];
      mem[10'd374] <= in[12223:12192];
      mem[10'd375] <= in[12191:12160];
      mem[10'd376] <= in[12159:12128];
      mem[10'd377] <= in[12127:12096];
      mem[10'd378] <= in[12095:12064];
      mem[10'd379] <= in[12063:12032];
      mem[10'd380] <= in[12031:12000];
      mem[10'd381] <= in[11999:11968];
      mem[10'd382] <= in[11967:11936];
      mem[10'd383] <= in[11935:11904];
      mem[10'd384] <= in[11903:11872];
      mem[10'd385] <= in[11871:11840];
      mem[10'd386] <= in[11839:11808];
      mem[10'd387] <= in[11807:11776];
      mem[10'd388] <= in[11775:11744];
      mem[10'd389] <= in[11743:11712];
      mem[10'd390] <= in[11711:11680];
      mem[10'd391] <= in[11679:11648];
      mem[10'd392] <= in[11647:11616];
      mem[10'd393] <= in[11615:11584];
      mem[10'd394] <= in[11583:11552];
      mem[10'd395] <= in[11551:11520];
      mem[10'd396] <= in[11519:11488];
      mem[10'd397] <= in[11487:11456];
      mem[10'd398] <= in[11455:11424];
      mem[10'd399] <= in[11423:11392];
      mem[10'd400] <= in[11391:11360];
      mem[10'd401] <= in[11359:11328];
      mem[10'd402] <= in[11327:11296];
      mem[10'd403] <= in[11295:11264];
      mem[10'd404] <= in[11263:11232];
      mem[10'd405] <= in[11231:11200];
      mem[10'd406] <= in[11199:11168];
      mem[10'd407] <= in[11167:11136];
      mem[10'd408] <= in[11135:11104];
      mem[10'd409] <= in[11103:11072];
      mem[10'd410] <= in[11071:11040];
      mem[10'd411] <= in[11039:11008];
      mem[10'd412] <= in[11007:10976];
      mem[10'd413] <= in[10975:10944];
      mem[10'd414] <= in[10943:10912];
      mem[10'd415] <= in[10911:10880];
      mem[10'd416] <= in[10879:10848];
      mem[10'd417] <= in[10847:10816];
      mem[10'd418] <= in[10815:10784];
      mem[10'd419] <= in[10783:10752];
      mem[10'd420] <= in[10751:10720];
      mem[10'd421] <= in[10719:10688];
      mem[10'd422] <= in[10687:10656];
      mem[10'd423] <= in[10655:10624];
      mem[10'd424] <= in[10623:10592];
      mem[10'd425] <= in[10591:10560];
      mem[10'd426] <= in[10559:10528];
      mem[10'd427] <= in[10527:10496];
      mem[10'd428] <= in[10495:10464];
      mem[10'd429] <= in[10463:10432];
      mem[10'd430] <= in[10431:10400];
      mem[10'd431] <= in[10399:10368];
      mem[10'd432] <= in[10367:10336];
      mem[10'd433] <= in[10335:10304];
      mem[10'd434] <= in[10303:10272];
      mem[10'd435] <= in[10271:10240];
      mem[10'd436] <= in[10239:10208];
      mem[10'd437] <= in[10207:10176];
      mem[10'd438] <= in[10175:10144];
      mem[10'd439] <= in[10143:10112];
      mem[10'd440] <= in[10111:10080];
      mem[10'd441] <= in[10079:10048];
      mem[10'd442] <= in[10047:10016];
      mem[10'd443] <= in[10015:9984];
      mem[10'd444] <= in[9983:9952];
      mem[10'd445] <= in[9951:9920];
      mem[10'd446] <= in[9919:9888];
      mem[10'd447] <= in[9887:9856];
      mem[10'd448] <= in[9855:9824];
      mem[10'd449] <= in[9823:9792];
      mem[10'd450] <= in[9791:9760];
      mem[10'd451] <= in[9759:9728];
      mem[10'd452] <= in[9727:9696];
      mem[10'd453] <= in[9695:9664];
      mem[10'd454] <= in[9663:9632];
      mem[10'd455] <= in[9631:9600];
      mem[10'd456] <= in[9599:9568];
      mem[10'd457] <= in[9567:9536];
      mem[10'd458] <= in[9535:9504];
      mem[10'd459] <= in[9503:9472];
      mem[10'd460] <= in[9471:9440];
      mem[10'd461] <= in[9439:9408];
      mem[10'd462] <= in[9407:9376];
      mem[10'd463] <= in[9375:9344];
      mem[10'd464] <= in[9343:9312];
      mem[10'd465] <= in[9311:9280];
      mem[10'd466] <= in[9279:9248];
      mem[10'd467] <= in[9247:9216];
      mem[10'd468] <= in[9215:9184];
      mem[10'd469] <= in[9183:9152];
      mem[10'd470] <= in[9151:9120];
      mem[10'd471] <= in[9119:9088];
      mem[10'd472] <= in[9087:9056];
      mem[10'd473] <= in[9055:9024];
      mem[10'd474] <= in[9023:8992];
      mem[10'd475] <= in[8991:8960];
      mem[10'd476] <= in[8959:8928];
      mem[10'd477] <= in[8927:8896];
      mem[10'd478] <= in[8895:8864];
      mem[10'd479] <= in[8863:8832];
      mem[10'd480] <= in[8831:8800];
      mem[10'd481] <= in[8799:8768];
      mem[10'd482] <= in[8767:8736];
      mem[10'd483] <= in[8735:8704];
      mem[10'd484] <= in[8703:8672];
      mem[10'd485] <= in[8671:8640];
      mem[10'd486] <= in[8639:8608];
      mem[10'd487] <= in[8607:8576];
      mem[10'd488] <= in[8575:8544];
      mem[10'd489] <= in[8543:8512];
      mem[10'd490] <= in[8511:8480];
      mem[10'd491] <= in[8479:8448];
      mem[10'd492] <= in[8447:8416];
      mem[10'd493] <= in[8415:8384];
      mem[10'd494] <= in[8383:8352];
      mem[10'd495] <= in[8351:8320];
      mem[10'd496] <= in[8319:8288];
      mem[10'd497] <= in[8287:8256];
      mem[10'd498] <= in[8255:8224];
      mem[10'd499] <= in[8223:8192];
      mem[10'd500] <= in[8191:8160];
      mem[10'd501] <= in[8159:8128];
      mem[10'd502] <= in[8127:8096];
      mem[10'd503] <= in[8095:8064];
      mem[10'd504] <= in[8063:8032];
      mem[10'd505] <= in[8031:8000];
      mem[10'd506] <= in[7999:7968];
      mem[10'd507] <= in[7967:7936];
      mem[10'd508] <= in[7935:7904];
      mem[10'd509] <= in[7903:7872];
      mem[10'd510] <= in[7871:7840];
      mem[10'd511] <= in[7839:7808];
      mem[10'd512] <= in[7807:7776];
      mem[10'd513] <= in[7775:7744];
      mem[10'd514] <= in[7743:7712];
      mem[10'd515] <= in[7711:7680];
      mem[10'd516] <= in[7679:7648];
      mem[10'd517] <= in[7647:7616];
      mem[10'd518] <= in[7615:7584];
      mem[10'd519] <= in[7583:7552];
      mem[10'd520] <= in[7551:7520];
      mem[10'd521] <= in[7519:7488];
      mem[10'd522] <= in[7487:7456];
      mem[10'd523] <= in[7455:7424];
      mem[10'd524] <= in[7423:7392];
      mem[10'd525] <= in[7391:7360];
      mem[10'd526] <= in[7359:7328];
      mem[10'd527] <= in[7327:7296];
      mem[10'd528] <= in[7295:7264];
      mem[10'd529] <= in[7263:7232];
      mem[10'd530] <= in[7231:7200];
      mem[10'd531] <= in[7199:7168];
      mem[10'd532] <= in[7167:7136];
      mem[10'd533] <= in[7135:7104];
      mem[10'd534] <= in[7103:7072];
      mem[10'd535] <= in[7071:7040];
      mem[10'd536] <= in[7039:7008];
      mem[10'd537] <= in[7007:6976];
      mem[10'd538] <= in[6975:6944];
      mem[10'd539] <= in[6943:6912];
      mem[10'd540] <= in[6911:6880];
      mem[10'd541] <= in[6879:6848];
      mem[10'd542] <= in[6847:6816];
      mem[10'd543] <= in[6815:6784];
      mem[10'd544] <= in[6783:6752];
      mem[10'd545] <= in[6751:6720];
      mem[10'd546] <= in[6719:6688];
      mem[10'd547] <= in[6687:6656];
      mem[10'd548] <= in[6655:6624];
      mem[10'd549] <= in[6623:6592];
      mem[10'd550] <= in[6591:6560];
      mem[10'd551] <= in[6559:6528];
      mem[10'd552] <= in[6527:6496];
      mem[10'd553] <= in[6495:6464];
      mem[10'd554] <= in[6463:6432];
      mem[10'd555] <= in[6431:6400];
      mem[10'd556] <= in[6399:6368];
      mem[10'd557] <= in[6367:6336];
      mem[10'd558] <= in[6335:6304];
      mem[10'd559] <= in[6303:6272];
      mem[10'd560] <= in[6271:6240];
      mem[10'd561] <= in[6239:6208];
      mem[10'd562] <= in[6207:6176];
      mem[10'd563] <= in[6175:6144];
      mem[10'd564] <= in[6143:6112];
      mem[10'd565] <= in[6111:6080];
      mem[10'd566] <= in[6079:6048];
      mem[10'd567] <= in[6047:6016];
      mem[10'd568] <= in[6015:5984];
      mem[10'd569] <= in[5983:5952];
      mem[10'd570] <= in[5951:5920];
      mem[10'd571] <= in[5919:5888];
      mem[10'd572] <= in[5887:5856];
      mem[10'd573] <= in[5855:5824];
      mem[10'd574] <= in[5823:5792];
      mem[10'd575] <= in[5791:5760];
      mem[10'd576] <= in[5759:5728];
      mem[10'd577] <= in[5727:5696];
      mem[10'd578] <= in[5695:5664];
      mem[10'd579] <= in[5663:5632];
      mem[10'd580] <= in[5631:5600];
      mem[10'd581] <= in[5599:5568];
      mem[10'd582] <= in[5567:5536];
      mem[10'd583] <= in[5535:5504];
      mem[10'd584] <= in[5503:5472];
      mem[10'd585] <= in[5471:5440];
      mem[10'd586] <= in[5439:5408];
      mem[10'd587] <= in[5407:5376];
      mem[10'd588] <= in[5375:5344];
      mem[10'd589] <= in[5343:5312];
      mem[10'd590] <= in[5311:5280];
      mem[10'd591] <= in[5279:5248];
      mem[10'd592] <= in[5247:5216];
      mem[10'd593] <= in[5215:5184];
      mem[10'd594] <= in[5183:5152];
      mem[10'd595] <= in[5151:5120];
      mem[10'd596] <= in[5119:5088];
      mem[10'd597] <= in[5087:5056];
      mem[10'd598] <= in[5055:5024];
      mem[10'd599] <= in[5023:4992];
      mem[10'd600] <= in[4991:4960];
      mem[10'd601] <= in[4959:4928];
      mem[10'd602] <= in[4927:4896];
      mem[10'd603] <= in[4895:4864];
      mem[10'd604] <= in[4863:4832];
      mem[10'd605] <= in[4831:4800];
      mem[10'd606] <= in[4799:4768];
      mem[10'd607] <= in[4767:4736];
      mem[10'd608] <= in[4735:4704];
      mem[10'd609] <= in[4703:4672];
      mem[10'd610] <= in[4671:4640];
      mem[10'd611] <= in[4639:4608];
      mem[10'd612] <= in[4607:4576];
      mem[10'd613] <= in[4575:4544];
      mem[10'd614] <= in[4543:4512];
      mem[10'd615] <= in[4511:4480];
      mem[10'd616] <= in[4479:4448];
      mem[10'd617] <= in[4447:4416];
      mem[10'd618] <= in[4415:4384];
      mem[10'd619] <= in[4383:4352];
      mem[10'd620] <= in[4351:4320];
      mem[10'd621] <= in[4319:4288];
      mem[10'd622] <= in[4287:4256];
      mem[10'd623] <= in[4255:4224];
      mem[10'd624] <= in[4223:4192];
      mem[10'd625] <= in[4191:4160];
      mem[10'd626] <= in[4159:4128];
      mem[10'd627] <= in[4127:4096];
      mem[10'd628] <= in[4095:4064];
      mem[10'd629] <= in[4063:4032];
      mem[10'd630] <= in[4031:4000];
      mem[10'd631] <= in[3999:3968];
      mem[10'd632] <= in[3967:3936];
      mem[10'd633] <= in[3935:3904];
      mem[10'd634] <= in[3903:3872];
      mem[10'd635] <= in[3871:3840];
      mem[10'd636] <= in[3839:3808];
      mem[10'd637] <= in[3807:3776];
      mem[10'd638] <= in[3775:3744];
      mem[10'd639] <= in[3743:3712];
      mem[10'd640] <= in[3711:3680];
      mem[10'd641] <= in[3679:3648];
      mem[10'd642] <= in[3647:3616];
      mem[10'd643] <= in[3615:3584];
      mem[10'd644] <= in[3583:3552];
      mem[10'd645] <= in[3551:3520];
      mem[10'd646] <= in[3519:3488];
      mem[10'd647] <= in[3487:3456];
      mem[10'd648] <= in[3455:3424];
      mem[10'd649] <= in[3423:3392];
      mem[10'd650] <= in[3391:3360];
      mem[10'd651] <= in[3359:3328];
      mem[10'd652] <= in[3327:3296];
      mem[10'd653] <= in[3295:3264];
      mem[10'd654] <= in[3263:3232];
      mem[10'd655] <= in[3231:3200];
      mem[10'd656] <= in[3199:3168];
      mem[10'd657] <= in[3167:3136];
      mem[10'd658] <= in[3135:3104];
      mem[10'd659] <= in[3103:3072];
      mem[10'd660] <= in[3071:3040];
      mem[10'd661] <= in[3039:3008];
      mem[10'd662] <= in[3007:2976];
      mem[10'd663] <= in[2975:2944];
      mem[10'd664] <= in[2943:2912];
      mem[10'd665] <= in[2911:2880];
      mem[10'd666] <= in[2879:2848];
      mem[10'd667] <= in[2847:2816];
      mem[10'd668] <= in[2815:2784];
      mem[10'd669] <= in[2783:2752];
      mem[10'd670] <= in[2751:2720];
      mem[10'd671] <= in[2719:2688];
      mem[10'd672] <= in[2687:2656];
      mem[10'd673] <= in[2655:2624];
      mem[10'd674] <= in[2623:2592];
      mem[10'd675] <= in[2591:2560];
      mem[10'd676] <= in[2559:2528];
      mem[10'd677] <= in[2527:2496];
      mem[10'd678] <= in[2495:2464];
      mem[10'd679] <= in[2463:2432];
      mem[10'd680] <= in[2431:2400];
      mem[10'd681] <= in[2399:2368];
      mem[10'd682] <= in[2367:2336];
      mem[10'd683] <= in[2335:2304];
      mem[10'd684] <= in[2303:2272];
      mem[10'd685] <= in[2271:2240];
      mem[10'd686] <= in[2239:2208];
      mem[10'd687] <= in[2207:2176];
      mem[10'd688] <= in[2175:2144];
      mem[10'd689] <= in[2143:2112];
      mem[10'd690] <= in[2111:2080];
      mem[10'd691] <= in[2079:2048];
      mem[10'd692] <= in[2047:2016];
      mem[10'd693] <= in[2015:1984];
      mem[10'd694] <= in[1983:1952];
      mem[10'd695] <= in[1951:1920];
      mem[10'd696] <= in[1919:1888];
      mem[10'd697] <= in[1887:1856];
      mem[10'd698] <= in[1855:1824];
      mem[10'd699] <= in[1823:1792];
      mem[10'd700] <= in[1791:1760];
      mem[10'd701] <= in[1759:1728];
      mem[10'd702] <= in[1727:1696];
      mem[10'd703] <= in[1695:1664];
      mem[10'd704] <= in[1663:1632];
      mem[10'd705] <= in[1631:1600];
      mem[10'd706] <= in[1599:1568];
      mem[10'd707] <= in[1567:1536];
      mem[10'd708] <= in[1535:1504];
      mem[10'd709] <= in[1503:1472];
      mem[10'd710] <= in[1471:1440];
      mem[10'd711] <= in[1439:1408];
      mem[10'd712] <= in[1407:1376];
      mem[10'd713] <= in[1375:1344];
      mem[10'd714] <= in[1343:1312];
      mem[10'd715] <= in[1311:1280];
      mem[10'd716] <= in[1279:1248];
      mem[10'd717] <= in[1247:1216];
      mem[10'd718] <= in[1215:1184];
      mem[10'd719] <= in[1183:1152];
      mem[10'd720] <= in[1151:1120];
      mem[10'd721] <= in[1119:1088];
      mem[10'd722] <= in[1087:1056];
      mem[10'd723] <= in[1055:1024];
      mem[10'd724] <= in[1023:992];
      mem[10'd725] <= in[991:960];
      mem[10'd726] <= in[959:928];
      mem[10'd727] <= in[927:896];
      mem[10'd728] <= in[895:864];
      mem[10'd729] <= in[863:832];
      mem[10'd730] <= in[831:800];
      mem[10'd731] <= in[799:768];
      mem[10'd732] <= in[767:736];
      mem[10'd733] <= in[735:704];
      mem[10'd734] <= in[703:672];
      mem[10'd735] <= in[671:640];
      mem[10'd736] <= in[639:608];
      mem[10'd737] <= in[607:576];
      mem[10'd738] <= in[575:544];
      mem[10'd739] <= in[543:512];
      mem[10'd740] <= in[511:480];
      mem[10'd741] <= in[479:448];
      mem[10'd742] <= in[447:416];
      mem[10'd743] <= in[415:384];
      mem[10'd744] <= in[383:352];
      mem[10'd745] <= in[351:320];
      mem[10'd746] <= in[319:288];
      mem[10'd747] <= in[287:256];
      mem[10'd748] <= in[255:224];
      mem[10'd749] <= in[223:192];
      mem[10'd750] <= in[191:160];
      mem[10'd751] <= in[159:128];
      mem[10'd752] <= in[127:96];
      mem[10'd753] <= in[95:64];
      mem[10'd754] <= in[63:32];
      mem[10'd755] <= in[31:0];
    end
    if(w_en) begin
      data_out <= mem[r_addr];
	  //Increase move counter if move is non-zero
	  if(mem[r_addr] != 32'd00000) begin
		move_counter = move_counter + 1;
	  end
	  //Done when all addresses have been read
	  if(r_addr == 10'd0755) begin
		done = 1'b1;
		move_counter_out <= move_counter;
	  end
	  r_addr <= r_addr + 10'd0001;
	  
    
    end
  end

endmodule